package uvm_def;
  import rtl_pkg::*;

endpackage
